module full_adder_test1();

    reg a , b, c ;

    wire sum , carry ; 

    FullAdder f(sum , carry , a , b ,c ); 

    initial 
        begin
            $monitor($time ,"a=%b , b=%b , c=%b , carry=%b , sum=%b" , a,b,c,sum,carry); 
             a=0; b=0; c=0;  
            #10 a=0; b=0; c=1; 
            #10 a=0; b=1; c=0; 
            #10 a=0; b=1; c=1; 
            #10 a=1; b=0; c=0; 
            #10 a=1; b=0; c=1; 
            #10 a=1; b=1; c=0; 
            #10 a=1; b=1; c=1;  

            #10 $finish ;
        end

endmodule